 `timescale 1ns/10ps
 module forwarding_unit(
						exe_mem_write_reg,
						mem_wb_write_reg,
						exe_mem_rd_addr,
						mem_wb_rd_addr,
						rs1_addr,
						rs2_addr,
						
						rs1_exe_hazard,
						rs1_mem_hazard,
						rs2_exe_hazard,
						rs2_mem_hazard					
						);
						
parameter DATA_SIZE  =32;
always_comb
begin
	
end

endmodule